`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 17.08.2025 22:04:05
// Design Name: 
// Module Name: concurrent_non_blocking
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module concurrent_non_blocking;
  reg clk, a, b;

  always @(posedge clk) begin
    a <= b;
    b <= a;
  end
endmodule
